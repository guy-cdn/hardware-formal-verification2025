package allocator_pkg;
   typedef enum reg [1:0] {IDLE, AQUIRE, PROCESS, RETURN} fsm_t;
endpackage // elevator_pkg
